module sand_update(
	input logic clock,
	input logic reset,

	input logic [15:0] region,
	input logic [15:0] floor,

	output logic [15:0] new_region,
	output logic [15:0] new_floor
    );


endmodule
